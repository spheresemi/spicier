Current Source Example
* 10mA current source with parallel resistors
* Expected: V(1) = 5V (10mA * 500 ohms)

I1 0 1 10m
R1 1 0 1k
R2 1 0 1k

.end
