DC Sweep of Voltage Divider
V1 1 0 DC 10
R1 1 2 1k
R2 2 0 1k
.dc V1 0 10 2
.end
