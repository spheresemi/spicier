RC Low-Pass Filter
V1 1 0 DC 5
R1 1 2 1k
C1 2 0 1u
.ac dec 5 1 1e6
.end
