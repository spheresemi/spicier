Nested DC Sweep Example - Transistor Curves
* Two voltage sources swept to trace I-V curves
V1 1 0 10
V2 2 0 5
R1 1 2 1k
R2 2 0 2k
.DC V1 0 10 2 V2 0 5 1
.END
