Voltage Divider Example
* Simple voltage divider with 10V source
* Expected: V(1)=10V, V(2)=5V

V1 1 0 DC 10
R1 1 2 1k
R2 2 0 1k

.end
