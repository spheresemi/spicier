Inductor DC Test
* At DC, inductor is a short circuit
* V(2) should equal V(1)

V1 1 0 10
L1 1 2 1m
R1 2 0 100

.end
