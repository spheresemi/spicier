RC Circuit (DC Analysis)
* At DC, capacitor is open circuit
* All current flows through R2

V1 1 0 12
R1 1 2 1k
C1 2 0 10u
R2 2 0 10k

.end
